`define CONTROLLER_STATE_READY 		0
`define CONTROLLER_STATE_ASSESS 	1
`define CONTROLLER_STATE_EXECUTE 	2

`define CONTROLLER_STATE_LOAD_BLOCK_NUMBER	10
`define CONTROLLER_STATE_LOAD_REG_NUMBER	11
`define CONTROLLER_STATE_LOAD_DATA			12
`define CONTROLLER_STATE_LOAD_INSTR			13

`define COMMAND_WRITE_BLOCK_INSTR 	8'b10010000
`define COMMAND_WRITE_BLOCK_REG 	8'b11100000
`define COMMAND_UPDATE_BLOCK_REG 	8'b11100001
`define COMMAND_ALLOC_SRAM_DELAY 	8'b00100000

`define INSTR 		32'h1
`define DATA 		32'h2
`define REG_NO 		32'h3
`define BLOCK_NO 	32'h4
