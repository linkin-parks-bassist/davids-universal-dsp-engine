`define LUT_HANDLE_WIDTH 8

`define LUT_FRAC_WIDTH 4
