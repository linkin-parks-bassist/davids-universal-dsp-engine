`define CONTROLLER_STATE_READY 		0
`define CONTROLLER_STATE_ASSESS 	1
`define CONTROLLER_STATE_EXECUTE 	2
`define CONTROLLER_STATE_SWAP_PAUSE	3
`define CONTROLLER_STATE_SWAP_WAIT 	4
`define CONTROLLER_STATE_RESET_WAIT 5
`define CONTROLLER_STATE_PAUSE		6

`define CONTROLLER_STATE_BEGIN				6

`define CONTROLLER_STATE_LOAD_BLOCK_NUMBER	10
`define CONTROLLER_STATE_LOAD_REG_NUMBER	11
`define CONTROLLER_STATE_LOAD_DATA			12
`define CONTROLLER_STATE_LOAD_INSTR			13

`define CONTROLLER_STATE_GET_BLOCK_NUMBER	10
`define CONTROLLER_STATE_GET_REG_NUMBER		11
`define CONTROLLER_STATE_GET_DATA			12
`define CONTROLLER_STATE_GET_INSTR			13
`define CONTROLLER_STATE_GET_DELAY			23

`define CONTROLLER_STATE_WRITE_BLOCK_INSTR 		14
`define CONTROLLER_STATE_WRITE_BLOCK_REG 		15
`define CONTROLLER_STATE_WRITE_BLOCK_REG_WAIT 	16
`define CONTROLLER_STATE_UPDATE_BLOCK_REG 		17
`define CONTROLLER_STATE_ALLOC_SRAM_DELAY 		18
`define CONTROLLER_STATE_SWAP_PIPELINES 		19
`define CONTROLLER_STATE_RESET_PIPELINE 		20
`define CONTROLLER_STATE_SET_INPUT_GAIN 		21
`define CONTROLLER_STATE_SET_OUTPUT_GAIN 		22
`define CONTROLLER_STATE_COMMIT_REG_UPDATES		23

`define COMMAND_WRITE_BLOCK_INSTR 	8'b10010000
`define COMMAND_WRITE_BLOCK_REG 	8'b11100000
`define COMMAND_UPDATE_BLOCK_REG 	8'b11101000
`define COMMAND_ALLOC_SRAM_DELAY 	8'b00100000
`define COMMAND_SWAP_PIPELINES 		8'b00000001
`define COMMAND_RESET_PIPELINE 		8'b00001001
`define COMMAND_SET_INPUT_GAIN 		8'b00000010
`define COMMAND_SET_OUTPUT_GAIN 	8'b00000011
`define COMMAND_COMMIT_REG_UPDATES 	8'b00001010

`define INSTR 		32'h1
`define DATA 		32'h2
`define REG_NO 		32'h3
`define BLOCK_NO 	32'h4
