`define CORE_STATE_READY 				0
`define CORE_STATE_BLOCK_START			1
`define CORE_STATE_FETCH_SRC_A			2
`define CORE_STATE_FETCH_SRC_A_2		3
`define CORE_STATE_FETCH_SRC_B			5
`define CORE_STATE_FETCH_SRC_B_2		6
`define CORE_STATE_FETCH_SRC_C			7
`define CORE_STATE_FETCH_SRC_C_2		8
`define CORE_STATE_FINISH_BLOCK			10
`define CORE_STATE_CONTINUE				11
`define CORE_STATE_DISPATCH				12
`define CORE_STATE_FINISH				13
`define CORE_STATE_COMMAND				14

`define CORE_STATE_ADD_1 			0110
`define CORE_STATE_ADD_2 			0210
`define CORE_STATE_SUB_1 			0120
`define CORE_STATE_SUB_2 			0220
`define CORE_STATE_MUL_1 			0160
`define CORE_STATE_MUL_2 			0260
`define CORE_STATE_MUL_3 			0360
`define CORE_STATE_MUL_4 			0460
`define CORE_STATE_MAD_1			0170
`define CORE_STATE_MAD_2			0270
`define CORE_STATE_MAD_3			0370
`define CORE_STATE_MAD_4			0470
`define CORE_STATE_MAD_5			0570
`define CORE_STATE_MAD_6			0670
`define CORE_STATE_LUT_1			0190
`define CORE_STATE_LUT_2			0290
`define CORE_STATE_LUT_3			0390
`define CORE_STATE_ENVD_1 			1100
`define CORE_STATE_DELAY_READ_1 	1110
`define CORE_STATE_DELAY_READ_2 	2110
`define CORE_STATE_DELAY_READ_3 	3110
`define CORE_STATE_DELAY_READ_4 	4110
`define CORE_STATE_DELAY_READ_5 	5110
`define CORE_STATE_DELAY_READ_6 	6110
`define CORE_STATE_DELAY_WRITE_1 	1120
`define CORE_STATE_DELAY_WRITE_2 	2120
`define CORE_STATE_DELAY_WRITE_3 	3120
`define CORE_STATE_DELAY_WRITE_4 	4120
`define CORE_STATE_DELAY_WRITE_5 	5120
`define CORE_STATE_DELAY_WRITE_6 	6120
`define CORE_STATE_SAVE_1 			1130
`define CORE_STATE_SAVE_2 			2130
`define CORE_STATE_LOAD_1			1140
`define CORE_STATE_MOV_1 			1150
`define CORE_STATE_CLAMP_1 			1160
`define CORE_STATE_MAC_1			1180
`define CORE_STATE_MAC_2			2180
`define CORE_STATE_MAC_3			3180
`define CORE_STATE_MAC_4			4180
`define CORE_STATE_MAC_5			5180
`define CORE_STATE_MAC_6			6180
